*** SPICE deck for cell NAND{ic} from library NAND
*** Created on Wed Aug 03, 2022 02:18:29
*** Last revised on Tue Aug 09, 2022 02:08:48
*** Written on Tue Aug 09, 2022 02:08:51 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: NAND{ic}

* Spice Code nodes in cell cell 'NAND{ic}'
vdd vdd 0 dc 1.8
va A 0 pulse (0 1.8 0 1n 1n 10n 20n)
vb B 0 pulse (0 1.8 0 1n 1n 20n 40n)
.tran 1n 100n
.include C:\Users\Mahmud Suhaimi\Desktop\EDA-Tool-1\tsmc_018um_model.txt
.END
